// The classic. Run with `v run helloworld.v`
module main

fn main() {
	println('Hello World, Hello V!')
}
